module andgate(y,a,b);
output y;
input a,b;
and a1(y,a,b);
endmodule