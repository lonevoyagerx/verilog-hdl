module encoder_tb;
reg[3:0] d;
wire[1:0]y;

encoder uut(d,y);

initial begin
    $dumpfile("encoder.vcd");
    $dumpvars(0,encoder_tb);
    $monitor("d=%b y=%b",d,y);

    d = 4'b0001;#10;
    d = 4'b0010;#10;
    d = 4'b0100;#10;
    d = 4'b1000;#10;

    $finish;
end
endmodule
