module orgate(y,a,b);
output y;
input a,b;
or a1(y,a,b);
endmodule