module xorgate(y,a,b);
output y;
input a,b;
xor a1(y,a,b);
endmodule