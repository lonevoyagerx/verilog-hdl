module norgate(y,a,b);
output y;
input a,b;
nor a1(y,a,b);
endmodule