module xnorgate(y,a,b);
output y;
input a,b;
xnor a1(y,a,b);
endmodule