module not_gate(a,y);
input a;
output y;
not a1(y,a);
endmodule