module full_sub_tb;
reg a,b,bin;
wire diff,borr;
full_sub uut (.diff(diff), .borr(borr), .a(a), .b(b), .bin(bin));

initial begin
    $dumpfile("dump.vcd");
    $dumpvars(0,full_sub_tb);
    $monitor("a = %b b = %b bin = %b diff = %b borr = %b",a,b,bin,diff,borr);

    a=0; b=0; bin=0; #10;
    a=0; b=0; bin=1; #10;
    a=0; b=1; bin=0; #10;
    a=0; b=1; bin=1; #10;
    a=1; b=0; bin=0; #10;
    a=1; b=0; bin=1; #10;
    a=1; b=1; bin=0; #10;
    a=1; b=1; bin=1; #10;

    $finish;
end
endmodule